module Processador();

endmodule